module top_module (
    output out);
    assign out = 0;
endmodule
